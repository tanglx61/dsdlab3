library verilog;
use verilog.vl_types.all;
entity g58_lab3_vlg_vec_tst is
end g58_lab3_vlg_vec_tst;

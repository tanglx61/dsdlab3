-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Wed Mar 15 14:29:01 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY g58_stack52 IS 
	PORT
	(
		enable :  IN  STD_LOGIC;
		rst :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		addr :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		data :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		mode :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		empty :  OUT  STD_LOGIC;
		full :  OUT  STD_LOGIC;
		num :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		value :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END g58_stack52;

ARCHITECTURE bdf_type OF g58_stack52 IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT lpm_ff_0
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_0: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_0: COMPONENT IS true;

COMPONENT lpm_ff_10
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_10: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_10: COMPONENT IS true;

COMPONENT lpm_ff_100
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_100: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_100: COMPONENT IS true;

COMPONENT lpm_ff_101
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_101: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_101: COMPONENT IS true;

COMPONENT lpm_ff_104
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_104: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_104: COMPONENT IS true;

COMPONENT lpm_ff_105
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_105: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_105: COMPONENT IS true;

COMPONENT lpm_ff_12
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_12: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_12: COMPONENT IS true;

COMPONENT lpm_ff_16
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_16: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_16: COMPONENT IS true;

COMPONENT lpm_ff_17
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_17: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_17: COMPONENT IS true;

COMPONENT lpm_ff_18
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_18: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_18: COMPONENT IS true;

COMPONENT lpm_ff_2
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_2: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_2: COMPONENT IS true;

COMPONENT lpm_ff_20
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_20: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_20: COMPONENT IS true;

COMPONENT lpm_ff_28
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_28: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_28: COMPONENT IS true;

COMPONENT lpm_ff_30
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_30: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_30: COMPONENT IS true;

COMPONENT lpm_ff_31
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_31: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_31: COMPONENT IS true;

COMPONENT lpm_ff_32
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_32: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_32: COMPONENT IS true;

COMPONENT lpm_ff_33
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_33: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_33: COMPONENT IS true;

COMPONENT lpm_ff_34
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_34: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_34: COMPONENT IS true;

COMPONENT lpm_ff_35
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_35: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_35: COMPONENT IS true;

COMPONENT lpm_ff_38
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_38: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_38: COMPONENT IS true;

COMPONENT lpm_ff_39
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_39: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_39: COMPONENT IS true;

COMPONENT lpm_ff_40
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_40: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_40: COMPONENT IS true;

COMPONENT lpm_ff_42
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_42: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_42: COMPONENT IS true;

COMPONENT lpm_ff_50
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_50: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_50: COMPONENT IS true;

COMPONENT lpm_ff_52
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_52: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_52: COMPONENT IS true;

COMPONENT lpm_ff_53
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_53: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_53: COMPONENT IS true;

COMPONENT lpm_ff_54
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_54: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_54: COMPONENT IS true;

COMPONENT lpm_ff_55
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_55: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_55: COMPONENT IS true;

COMPONENT lpm_ff_56
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_56: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_56: COMPONENT IS true;

COMPONENT lpm_ff_57
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_57: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_57: COMPONENT IS true;

COMPONENT lpm_ff_60
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_60: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_60: COMPONENT IS true;

COMPONENT lpm_ff_61
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_61: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_61: COMPONENT IS true;

COMPONENT lpm_ff_62
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_62: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_62: COMPONENT IS true;

COMPONENT lpm_ff_7
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_7: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_7: COMPONENT IS true;

COMPONENT lpm_ff_74
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_74: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_74: COMPONENT IS true;

COMPONENT lpm_ff_75
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_75: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_75: COMPONENT IS true;

COMPONENT lpm_ff_76
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_76: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_76: COMPONENT IS true;

COMPONENT lpm_ff_77
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_77: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_77: COMPONENT IS true;

COMPONENT lpm_ff_78
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_78: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_78: COMPONENT IS true;

COMPONENT lpm_ff_79
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_79: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_79: COMPONENT IS true;

COMPONENT lpm_ff_8
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_8: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_8: COMPONENT IS true;

COMPONENT lpm_ff_80
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_80: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_80: COMPONENT IS true;

COMPONENT lpm_ff_81
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_81: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_81: COMPONENT IS true;

COMPONENT lpm_ff_82
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_82: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_82: COMPONENT IS true;

COMPONENT lpm_ff_83
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_83: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_83: COMPONENT IS true;

COMPONENT lpm_ff_84
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_84: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_84: COMPONENT IS true;

COMPONENT lpm_ff_86
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_86: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_86: COMPONENT IS true;

COMPONENT lpm_ff_9
	PORT(clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_9: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_9: COMPONENT IS true;

COMPONENT lpm_ff_94
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_94: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_94: COMPONENT IS true;

COMPONENT lpm_ff_96
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_96: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_96: COMPONENT IS true;

COMPONENT lpm_ff_97
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_97: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_97: COMPONENT IS true;

COMPONENT lpm_ff_98
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_98: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_98: COMPONENT IS true;

COMPONENT lpm_ff_99
	PORT(aclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_99: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_99: COMPONENT IS true;

TYPE ARRAY2D0 IS ARRAY (51 DOWNTO 0,5 DOWNTO 0) OF STD_LOGIC;

COMPONENT lpm_mux_5
	PORT(data : IN ARRAY2D0;
		 sel : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_mux_5: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_mux_5: COMPONENT IS true;

COMPONENT busmux_1
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_1: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_1: COMPONENT IS true;

COMPONENT busmux_102
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_102: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_102: COMPONENT IS true;

COMPONENT busmux_103
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_103: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_103: COMPONENT IS true;

COMPONENT busmux_11
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_11: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_11: COMPONENT IS true;

COMPONENT busmux_13
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_13: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_13: COMPONENT IS true;

COMPONENT busmux_14
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_14: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_14: COMPONENT IS true;

COMPONENT busmux_15
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_15: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_15: COMPONENT IS true;

COMPONENT busmux_19
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_19: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_19: COMPONENT IS true;

COMPONENT busmux_21
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_21: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_21: COMPONENT IS true;

COMPONENT busmux_22
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_22: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_22: COMPONENT IS true;

COMPONENT busmux_23
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_23: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_23: COMPONENT IS true;

COMPONENT busmux_24
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_24: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_24: COMPONENT IS true;

COMPONENT busmux_25
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_25: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_25: COMPONENT IS true;

COMPONENT busmux_26
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_26: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_26: COMPONENT IS true;

COMPONENT busmux_27
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_27: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_27: COMPONENT IS true;

COMPONENT busmux_29
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_29: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_29: COMPONENT IS true;

COMPONENT busmux_3
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_3: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_3: COMPONENT IS true;

COMPONENT busmux_36
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_36: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_36: COMPONENT IS true;

COMPONENT busmux_37
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_37: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_37: COMPONENT IS true;

COMPONENT busmux_4
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_4: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_4: COMPONENT IS true;

COMPONENT busmux_41
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_41: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_41: COMPONENT IS true;

COMPONENT busmux_43
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_43: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_43: COMPONENT IS true;

COMPONENT busmux_44
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_44: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_44: COMPONENT IS true;

COMPONENT busmux_45
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_45: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_45: COMPONENT IS true;

COMPONENT busmux_46
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_46: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_46: COMPONENT IS true;

COMPONENT busmux_47
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_47: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_47: COMPONENT IS true;

COMPONENT busmux_48
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_48: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_48: COMPONENT IS true;

COMPONENT busmux_49
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_49: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_49: COMPONENT IS true;

COMPONENT busmux_51
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_51: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_51: COMPONENT IS true;

COMPONENT busmux_58
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_58: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_58: COMPONENT IS true;

COMPONENT busmux_59
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_59: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_59: COMPONENT IS true;

COMPONENT busmux_6
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_6: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_6: COMPONENT IS true;

COMPONENT busmux_63
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_63: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_63: COMPONENT IS true;

COMPONENT busmux_64
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_64: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_64: COMPONENT IS true;

COMPONENT busmux_65
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_65: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_65: COMPONENT IS true;

COMPONENT busmux_66
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_66: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_66: COMPONENT IS true;

COMPONENT busmux_67
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_67: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_67: COMPONENT IS true;

COMPONENT busmux_68
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_68: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_68: COMPONENT IS true;

COMPONENT busmux_69
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_69: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_69: COMPONENT IS true;

COMPONENT busmux_70
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_70: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_70: COMPONENT IS true;

COMPONENT busmux_71
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_71: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_71: COMPONENT IS true;

COMPONENT busmux_72
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_72: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_72: COMPONENT IS true;

COMPONENT busmux_73
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_73: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_73: COMPONENT IS true;

COMPONENT busmux_85
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_85: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_85: COMPONENT IS true;

COMPONENT busmux_87
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_87: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_87: COMPONENT IS true;

COMPONENT busmux_88
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_88: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_88: COMPONENT IS true;

COMPONENT busmux_89
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_89: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_89: COMPONENT IS true;

COMPONENT busmux_90
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_90: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_90: COMPONENT IS true;

COMPONENT busmux_91
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_91: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_91: COMPONENT IS true;

COMPONENT busmux_92
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_92: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_92: COMPONENT IS true;

COMPONENT busmux_93
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_93: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_93: COMPONENT IS true;

COMPONENT busmux_95
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_95: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_95: COMPONENT IS true;

COMPONENT g58_pop_enable
	PORT(CLK : IN STD_LOGIC;
		 N : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 P_EN : OUT STD_LOGIC_VECTOR(51 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	a :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	aa :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	b :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	bb :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	c :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	cc :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	d :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	dd :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	e :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	ee :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	f :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	ff :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	g :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	gg :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	h :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	hh :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	i :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	ii :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	init :  STD_LOGIC;
SIGNAL	j :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	jj :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	k :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	kk :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	l :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	ll :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	m :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	mm :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	n :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	nn :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	o :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	oo :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	p :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	P_EN :  STD_LOGIC_VECTOR(51 DOWNTO 0);
SIGNAL	pp :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	q :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	qq :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	r :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	rr :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	s :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	sh :  STD_LOGIC;
SIGNAL	ss :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	t :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	tt :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	u :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	uu :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	v :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	vv :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	w :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	ww :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	x :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	xx :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	y :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	yy :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	z :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	zz :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC_VECTOR(5 DOWNTO 0);

SIGNAL	GDFX_TEMP_SIGNAL_0 :  ARRAY2D0;

BEGIN 

GDFX_TEMP_SIGNAL_0 <= (a(5 DOWNTO 0) & b(5 DOWNTO 0) & c(5 DOWNTO 0) & d(5 DOWNTO 0) & e(5 DOWNTO 0) & f(5 DOWNTO 0) & g(5 DOWNTO 0) & h(5 DOWNTO 0) & i(5 DOWNTO 0) & j(5 DOWNTO 0) & k(5 DOWNTO 0) & l(5 DOWNTO 0) & m(5 DOWNTO 0) & n(5 DOWNTO 0) & o(5 DOWNTO 0) & p(5 DOWNTO 0) & q(5 DOWNTO 0) & r(5 DOWNTO 0) & s(5 DOWNTO 0) & t(5 DOWNTO 0) & u(5 DOWNTO 0) & v(5 DOWNTO 0) & w(5 DOWNTO 0) & x(5 DOWNTO 0) & y(5 DOWNTO 0) & z(5 DOWNTO 0) & aa(5 DOWNTO 0) & bb(5 DOWNTO 0) & cc(5 DOWNTO 0) & dd(5 DOWNTO 0) & ee(5 DOWNTO 0) & ff(5 DOWNTO 0) & gg(5 DOWNTO 0) & hh(5 DOWNTO 0) & ii(5 DOWNTO 0) & jj(5 DOWNTO 0) & kk(5 DOWNTO 0) & ll(5 DOWNTO 0) & mm(5 DOWNTO 0) & nn(5 DOWNTO 0) & oo(5 DOWNTO 0) & pp(5 DOWNTO 0) & qq(5 DOWNTO 0) & rr(5 DOWNTO 0) & ss(5 DOWNTO 0) & tt(5 DOWNTO 0) & uu(5 DOWNTO 0) & vv(5 DOWNTO 0) & ww(5 DOWNTO 0) & xx(5 DOWNTO 0) & yy(5 DOWNTO 0) & zz(5 DOWNTO 0));


b2v_inst : lpm_ff_0
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(0),
		 sset => init,
		 data => SYNTHESIZED_WIRE_0,
		 q => zz);


b2v_inst1 : busmux_1
PORT MAP(sel => sh,
		 dataa => data,
		 datab => yy,
		 result => SYNTHESIZED_WIRE_0);


b2v_inst10 : lpm_ff_2
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(5),
		 sset => init,
		 data => SYNTHESIZED_WIRE_1,
		 q => uu);


b2v_inst100 : busmux_3
PORT MAP(sel => sh,
		 dataa => c,
		 datab => a,
		 result => SYNTHESIZED_WIRE_4);


b2v_inst101 : busmux_4
PORT MAP(sel => sh,
		 dataa => b,
		 datab => SYNTHESIZED_WIRE_2,
		 result => SYNTHESIZED_WIRE_5);


b2v_inst102 : g58_pop_enable
PORT MAP(CLK => clk,
		 N => addr,
		 P_EN => P_EN);


b2v_inst103 : lpm_mux_5
PORT MAP(data => GDFX_TEMP_SIGNAL_0,
		 sel => addr,
		 result => value);


init <= SYNTHESIZED_WIRE_3 AND mode(1);


SYNTHESIZED_WIRE_3 <= NOT(mode(0));



sh <= mode(0) AND mode(1);


b2v_inst11 : busmux_6
PORT MAP(sel => sh,
		 dataa => vv,
		 datab => tt,
		 result => SYNTHESIZED_WIRE_1);


b2v_inst110 : lpm_ff_7
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(50),
		 sset => init,
		 data => SYNTHESIZED_WIRE_4,
		 q => b);


b2v_inst111 : lpm_ff_8
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(51),
		 sset => init,
		 data => SYNTHESIZED_WIRE_5,
		 q => a);


b2v_inst112 : lpm_ff_9
PORT MAP(clock => clk,
		 sset => init,
		 q => SYNTHESIZED_WIRE_2);


b2v_inst12 : lpm_ff_10
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(6),
		 sset => init,
		 data => SYNTHESIZED_WIRE_6,
		 q => tt);


b2v_inst13 : busmux_11
PORT MAP(sel => sh,
		 dataa => uu,
		 datab => ss,
		 result => SYNTHESIZED_WIRE_6);


b2v_inst14 : lpm_ff_12
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(7),
		 sset => init,
		 data => SYNTHESIZED_WIRE_7,
		 q => ss);


b2v_inst15 : busmux_13
PORT MAP(sel => sh,
		 dataa => tt,
		 datab => rr,
		 result => SYNTHESIZED_WIRE_7);


b2v_inst16 : busmux_14
PORT MAP(sel => sh,
		 dataa => ss,
		 datab => qq,
		 result => SYNTHESIZED_WIRE_8);


b2v_inst17 : busmux_15
PORT MAP(sel => sh,
		 dataa => rr,
		 datab => pp,
		 result => SYNTHESIZED_WIRE_9);


b2v_inst18 : lpm_ff_16
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(8),
		 sset => init,
		 data => SYNTHESIZED_WIRE_8,
		 q => rr);


b2v_inst19 : lpm_ff_17
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(9),
		 sset => init,
		 data => SYNTHESIZED_WIRE_9,
		 q => qq);


b2v_inst2 : lpm_ff_18
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(1),
		 sset => init,
		 data => SYNTHESIZED_WIRE_10,
		 q => yy);


b2v_inst20 : busmux_19
PORT MAP(sel => sh,
		 dataa => qq,
		 datab => oo,
		 result => SYNTHESIZED_WIRE_14);


b2v_inst21 : lpm_ff_20
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(11),
		 sset => init,
		 data => SYNTHESIZED_WIRE_11,
		 q => oo);


b2v_inst22 : busmux_21
PORT MAP(sel => sh,
		 dataa => pp,
		 datab => nn,
		 result => SYNTHESIZED_WIRE_11);


b2v_inst23 : busmux_22
PORT MAP(sel => sh,
		 dataa => oo,
		 datab => mm,
		 result => SYNTHESIZED_WIRE_12);


b2v_inst24 : busmux_23
PORT MAP(sel => sh,
		 dataa => nn,
		 datab => ll,
		 result => SYNTHESIZED_WIRE_13);


b2v_inst25 : busmux_24
PORT MAP(sel => sh,
		 dataa => mm,
		 datab => kk,
		 result => SYNTHESIZED_WIRE_15);


b2v_inst26 : busmux_25
PORT MAP(sel => sh,
		 dataa => ll,
		 datab => jj,
		 result => SYNTHESIZED_WIRE_16);


b2v_inst27 : busmux_26
PORT MAP(sel => sh,
		 dataa => kk,
		 datab => ii,
		 result => SYNTHESIZED_WIRE_17);


b2v_inst28 : busmux_27
PORT MAP(sel => sh,
		 dataa => jj,
		 datab => hh,
		 result => SYNTHESIZED_WIRE_18);


b2v_inst29 : lpm_ff_28
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(12),
		 sset => init,
		 data => SYNTHESIZED_WIRE_12,
		 q => nn);


b2v_inst3 : busmux_29
PORT MAP(sel => sh,
		 dataa => zz,
		 datab => xx,
		 result => SYNTHESIZED_WIRE_10);


b2v_inst30 : lpm_ff_30
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(13),
		 sset => init,
		 data => SYNTHESIZED_WIRE_13,
		 q => mm);


b2v_inst31 : lpm_ff_31
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(10),
		 sset => init,
		 data => SYNTHESIZED_WIRE_14,
		 q => pp);


b2v_inst32 : lpm_ff_32
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(14),
		 sset => init,
		 data => SYNTHESIZED_WIRE_15,
		 q => ll);


b2v_inst33 : lpm_ff_33
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(15),
		 sset => init,
		 data => SYNTHESIZED_WIRE_16,
		 q => kk);


b2v_inst34 : lpm_ff_34
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(16),
		 sset => init,
		 data => SYNTHESIZED_WIRE_17,
		 q => jj);


b2v_inst35 : lpm_ff_35
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(17),
		 sset => init,
		 data => SYNTHESIZED_WIRE_18,
		 q => ii);


b2v_inst36 : busmux_36
PORT MAP(sel => sh,
		 dataa => ii,
		 datab => gg,
		 result => SYNTHESIZED_WIRE_19);


b2v_inst37 : busmux_37
PORT MAP(sel => sh,
		 dataa => hh,
		 datab => ff,
		 result => SYNTHESIZED_WIRE_20);


b2v_inst38 : lpm_ff_38
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(18),
		 sset => init,
		 data => SYNTHESIZED_WIRE_19,
		 q => hh);


b2v_inst39 : lpm_ff_39
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(19),
		 sset => init,
		 data => SYNTHESIZED_WIRE_20,
		 q => gg);


b2v_inst4 : lpm_ff_40
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(2),
		 sset => init,
		 data => SYNTHESIZED_WIRE_21,
		 q => xx);


b2v_inst40 : busmux_41
PORT MAP(sel => sh,
		 dataa => gg,
		 datab => ee,
		 result => SYNTHESIZED_WIRE_23);


b2v_inst41 : lpm_ff_42
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(21),
		 sset => init,
		 data => SYNTHESIZED_WIRE_22,
		 q => ee);


b2v_inst42 : busmux_43
PORT MAP(sel => sh,
		 dataa => ff,
		 datab => dd,
		 result => SYNTHESIZED_WIRE_22);


b2v_inst43 : busmux_44
PORT MAP(sel => sh,
		 dataa => ee,
		 datab => cc,
		 result => SYNTHESIZED_WIRE_24);


b2v_inst44 : busmux_45
PORT MAP(sel => sh,
		 dataa => dd,
		 datab => bb,
		 result => SYNTHESIZED_WIRE_25);


b2v_inst45 : busmux_46
PORT MAP(sel => sh,
		 dataa => cc,
		 datab => aa,
		 result => SYNTHESIZED_WIRE_26);


b2v_inst46 : busmux_47
PORT MAP(sel => sh,
		 dataa => bb,
		 datab => z,
		 result => SYNTHESIZED_WIRE_27);


b2v_inst47 : busmux_48
PORT MAP(sel => sh,
		 dataa => aa,
		 datab => y,
		 result => SYNTHESIZED_WIRE_28);


b2v_inst48 : busmux_49
PORT MAP(sel => sh,
		 dataa => z,
		 datab => x,
		 result => SYNTHESIZED_WIRE_29);


b2v_inst49 : lpm_ff_50
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(20),
		 sset => init,
		 data => SYNTHESIZED_WIRE_23,
		 q => ff);


b2v_inst5 : busmux_51
PORT MAP(sel => sh,
		 dataa => yy,
		 datab => ww,
		 result => SYNTHESIZED_WIRE_21);


b2v_inst50 : lpm_ff_52
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(22),
		 sset => init,
		 data => SYNTHESIZED_WIRE_24,
		 q => dd);


b2v_inst51 : lpm_ff_53
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(23),
		 sset => init,
		 data => SYNTHESIZED_WIRE_25,
		 q => cc);


b2v_inst52 : lpm_ff_54
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(24),
		 sset => init,
		 data => SYNTHESIZED_WIRE_26,
		 q => bb);


b2v_inst53 : lpm_ff_55
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(25),
		 sset => init,
		 data => SYNTHESIZED_WIRE_27,
		 q => aa);


b2v_inst54 : lpm_ff_56
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(26),
		 sset => init,
		 data => SYNTHESIZED_WIRE_28,
		 q => z);


b2v_inst55 : lpm_ff_57
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(27),
		 sset => init,
		 data => SYNTHESIZED_WIRE_29,
		 q => y);


b2v_inst56 : busmux_58
PORT MAP(sel => sh,
		 dataa => y,
		 datab => w,
		 result => SYNTHESIZED_WIRE_30);


b2v_inst57 : busmux_59
PORT MAP(sel => sh,
		 dataa => x,
		 datab => v,
		 result => SYNTHESIZED_WIRE_31);


b2v_inst58 : lpm_ff_60
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(28),
		 sset => init,
		 data => SYNTHESIZED_WIRE_30,
		 q => x);


b2v_inst59 : lpm_ff_61
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(29),
		 sset => init,
		 data => SYNTHESIZED_WIRE_31,
		 q => w);


b2v_inst6 : lpm_ff_62
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(3),
		 sset => init,
		 data => SYNTHESIZED_WIRE_32,
		 q => ww);


b2v_inst60 : busmux_63
PORT MAP(sel => sh,
		 dataa => w,
		 datab => u,
		 result => SYNTHESIZED_WIRE_33);


b2v_inst61 : busmux_64
PORT MAP(sel => sh,
		 dataa => v,
		 datab => t,
		 result => SYNTHESIZED_WIRE_34);


b2v_inst62 : busmux_65
PORT MAP(sel => sh,
		 dataa => u,
		 datab => s,
		 result => SYNTHESIZED_WIRE_35);


b2v_inst63 : busmux_66
PORT MAP(sel => sh,
		 dataa => t,
		 datab => r,
		 result => SYNTHESIZED_WIRE_36);


b2v_inst64 : busmux_67
PORT MAP(sel => sh,
		 dataa => s,
		 datab => q,
		 result => SYNTHESIZED_WIRE_37);


b2v_inst65 : busmux_68
PORT MAP(sel => sh,
		 dataa => r,
		 datab => p,
		 result => SYNTHESIZED_WIRE_38);


b2v_inst66 : busmux_69
PORT MAP(sel => sh,
		 dataa => q,
		 datab => o,
		 result => SYNTHESIZED_WIRE_39);


b2v_inst67 : busmux_70
PORT MAP(sel => sh,
		 dataa => p,
		 datab => n,
		 result => SYNTHESIZED_WIRE_40);


b2v_inst68 : busmux_71
PORT MAP(sel => sh,
		 dataa => o,
		 datab => m,
		 result => SYNTHESIZED_WIRE_41);


b2v_inst69 : busmux_72
PORT MAP(sel => sh,
		 dataa => n,
		 datab => l,
		 result => SYNTHESIZED_WIRE_42);


b2v_inst7 : busmux_73
PORT MAP(sel => sh,
		 dataa => xx,
		 datab => vv,
		 result => SYNTHESIZED_WIRE_32);


b2v_inst70 : lpm_ff_74
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(30),
		 sset => init,
		 data => SYNTHESIZED_WIRE_33,
		 q => v);


b2v_inst71 : lpm_ff_75
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(31),
		 sset => init,
		 data => SYNTHESIZED_WIRE_34,
		 q => u);


b2v_inst72 : lpm_ff_76
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(32),
		 sset => init,
		 data => SYNTHESIZED_WIRE_35,
		 q => t);


b2v_inst73 : lpm_ff_77
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(33),
		 sset => init,
		 data => SYNTHESIZED_WIRE_36,
		 q => s);


b2v_inst74 : lpm_ff_78
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(34),
		 sset => init,
		 data => SYNTHESIZED_WIRE_37,
		 q => r);


b2v_inst75 : lpm_ff_79
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(35),
		 sset => init,
		 data => SYNTHESIZED_WIRE_38,
		 q => q);


b2v_inst76 : lpm_ff_80
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(36),
		 sset => init,
		 data => SYNTHESIZED_WIRE_39,
		 q => p);


b2v_inst77 : lpm_ff_81
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(37),
		 sset => init,
		 data => SYNTHESIZED_WIRE_40,
		 q => o);


b2v_inst78 : lpm_ff_82
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(38),
		 sset => init,
		 data => SYNTHESIZED_WIRE_41,
		 q => n);


b2v_inst79 : lpm_ff_83
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(39),
		 sset => init,
		 data => SYNTHESIZED_WIRE_42,
		 q => m);


b2v_inst8 : lpm_ff_84
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(4),
		 sset => init,
		 data => SYNTHESIZED_WIRE_43,
		 q => vv);


b2v_inst80 : busmux_85
PORT MAP(sel => sh,
		 dataa => m,
		 datab => k,
		 result => SYNTHESIZED_WIRE_45);


b2v_inst81 : lpm_ff_86
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(41),
		 sset => init,
		 data => SYNTHESIZED_WIRE_44,
		 q => k);


b2v_inst82 : busmux_87
PORT MAP(sel => sh,
		 dataa => l,
		 datab => j,
		 result => SYNTHESIZED_WIRE_44);


b2v_inst83 : busmux_88
PORT MAP(sel => sh,
		 dataa => k,
		 datab => i,
		 result => SYNTHESIZED_WIRE_46);


b2v_inst84 : busmux_89
PORT MAP(sel => sh,
		 dataa => j,
		 datab => h,
		 result => SYNTHESIZED_WIRE_47);


b2v_inst85 : busmux_90
PORT MAP(sel => sh,
		 dataa => i,
		 datab => g,
		 result => SYNTHESIZED_WIRE_48);


b2v_inst86 : busmux_91
PORT MAP(sel => sh,
		 dataa => h,
		 datab => f,
		 result => SYNTHESIZED_WIRE_49);


b2v_inst87 : busmux_92
PORT MAP(sel => sh,
		 dataa => g,
		 datab => e,
		 result => SYNTHESIZED_WIRE_50);


b2v_inst88 : busmux_93
PORT MAP(sel => sh,
		 dataa => f,
		 datab => d,
		 result => SYNTHESIZED_WIRE_51);


b2v_inst89 : lpm_ff_94
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(40),
		 sset => init,
		 data => SYNTHESIZED_WIRE_45,
		 q => l);


b2v_inst9 : busmux_95
PORT MAP(sel => sh,
		 dataa => ww,
		 datab => uu,
		 result => SYNTHESIZED_WIRE_43);


b2v_inst90 : lpm_ff_96
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(42),
		 sset => init,
		 data => SYNTHESIZED_WIRE_46,
		 q => j);


b2v_inst91 : lpm_ff_97
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(43),
		 sset => init,
		 data => SYNTHESIZED_WIRE_47,
		 q => i);


b2v_inst92 : lpm_ff_98
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(44),
		 sset => init,
		 data => SYNTHESIZED_WIRE_48,
		 q => h);


b2v_inst93 : lpm_ff_99
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(45),
		 sset => init,
		 data => SYNTHESIZED_WIRE_49,
		 q => g);


b2v_inst94 : lpm_ff_100
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(46),
		 sset => init,
		 data => SYNTHESIZED_WIRE_50,
		 q => f);


b2v_inst95 : lpm_ff_101
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(47),
		 sset => init,
		 data => SYNTHESIZED_WIRE_51,
		 q => e);


b2v_inst96 : busmux_102
PORT MAP(sel => sh,
		 dataa => e,
		 datab => c,
		 result => SYNTHESIZED_WIRE_52);


b2v_inst97 : busmux_103
PORT MAP(sel => sh,
		 dataa => d,
		 datab => b,
		 result => SYNTHESIZED_WIRE_53);


b2v_inst98 : lpm_ff_104
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(48),
		 sset => init,
		 data => SYNTHESIZED_WIRE_52,
		 q => d);


b2v_inst99 : lpm_ff_105
PORT MAP(aclr => rst,
		 clock => clk,
		 enable => P_EN(49),
		 sset => init,
		 data => SYNTHESIZED_WIRE_53,
		 q => c);


END bdf_type;
library verilog;
use verilog.vl_types.all;
entity g58_pulse_gen_test_vlg_vec_tst is
end g58_pulse_gen_test_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity g58_pulse_gen_test_vlg_check_tst is
    port(
        pulse           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g58_pulse_gen_test_vlg_check_tst;
